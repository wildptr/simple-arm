module asr(
  input [32:0] in,
  input [ 7:0] sh,
  output reg [32:0] out
);

always @* begin
  case (sh)
    8'd 0: out = in;
    8'd 1: out = {{ 1{in[32]}}, in[32: 1]};
    8'd 2: out = {{ 2{in[32]}}, in[32: 2]};
    8'd 3: out = {{ 3{in[32]}}, in[32: 3]};
    8'd 4: out = {{ 4{in[32]}}, in[32: 4]};
    8'd 5: out = {{ 5{in[32]}}, in[32: 5]};
    8'd 6: out = {{ 6{in[32]}}, in[32: 6]};
    8'd 7: out = {{ 7{in[32]}}, in[32: 7]};
    8'd 8: out = {{ 8{in[32]}}, in[32: 8]};
    8'd 9: out = {{ 9{in[32]}}, in[32: 9]};
    8'd10: out = {{10{in[32]}}, in[32:10]};
    8'd11: out = {{11{in[32]}}, in[32:11]};
    8'd12: out = {{12{in[32]}}, in[32:12]};
    8'd13: out = {{13{in[32]}}, in[32:13]};
    8'd14: out = {{14{in[32]}}, in[32:14]};
    8'd15: out = {{15{in[32]}}, in[32:15]};
    8'd16: out = {{16{in[32]}}, in[32:16]};
    8'd17: out = {{17{in[32]}}, in[32:17]};
    8'd18: out = {{18{in[32]}}, in[32:18]};
    8'd19: out = {{19{in[32]}}, in[32:19]};
    8'd20: out = {{20{in[32]}}, in[32:20]};
    8'd21: out = {{21{in[32]}}, in[32:21]};
    8'd22: out = {{22{in[32]}}, in[32:22]};
    8'd23: out = {{23{in[32]}}, in[32:23]};
    8'd24: out = {{24{in[32]}}, in[32:24]};
    8'd25: out = {{25{in[32]}}, in[32:25]};
    8'd26: out = {{26{in[32]}}, in[32:26]};
    8'd27: out = {{27{in[32]}}, in[32:27]};
    8'd28: out = {{28{in[32]}}, in[32:28]};
    8'd29: out = {{29{in[32]}}, in[32:29]};
    8'd30: out = {{30{in[32]}}, in[32:30]};
    8'd31: out = {{31{in[32]}}, in[32:31]};
    default: out = {33{in[32]}};
  endcase
end

endmodule
